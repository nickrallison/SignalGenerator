module data_loader #(ADDRESS_SIZE=8, DATA_SIZE=8, DATA_LEN=256) (
    input logic i_clk,
    input logic i_res,
    input logic i_data,
    output logic o_data
);



endmodule