module repeater #() (
    input logic i_clk,
    input logic i_res,
    input logic i_data,
    output logic o_data
);
